* /home/ganapathisubramanian28/Downloads/ganapathijohnsoncounter/johnsoncounter/johnsoncounter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 05 Mar 2022 06:28:12 AM UTC

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M4  Net-_M3-Pad1_ Net-_M1-Pad1_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M6  Net-_M1-Pad2_ Net-_M3-Pad1_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ GND GND mosfet_n		
M3  Net-_M3-Pad1_ Net-_M1-Pad1_ GND GND mosfet_n		
M5  Net-_M1-Pad2_ Net-_M3-Pad1_ GND GND mosfet_n		
U1  clk plot_v1		
v1  Net-_M2-Pad3_ GND DC		
U3  clk Net-_U3-Pad2_ Net-_U2-Pad1_ Net-_U2-Pad2_ adc_bridge_2		
U4  Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ o3 o2 o1 o0 dac_bridge_4		
U5  o3 plot_v1		
U6  o2 plot_v1		
U7  o1 plot_v1		
U8  o0 plot_v1		
v2  Net-_U3-Pad2_ GND pulse		
R1  Net-_M1-Pad2_ clk 10k		
R2  clk GND 10k		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ johnson		

.end
